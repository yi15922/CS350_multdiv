//module divControl(add, sub, shiftProductDiv, nop, )