module multdiv(
	data_operandA, data_operandB, 
	ctrl_MULT, ctrl_DIV, 
	clock, 
	data_result, data_exception, data_resultRDY);

    input [31:0] data_operandA, data_operandB;
    input ctrl_MULT, ctrl_DIV, clock;

    output [31:0] data_result;
    output data_exception, data_resultRDY;

    // add your code here

    wire shiftMultiplicand; 
    wire [31:0] multiplicand;
    assign multiplicand = shiftMultiplicand ? multiplicand << 1 : multiplicand; 

    //register64 reg()

endmodule