module div(data_operandA, data_operandB, ctrl_DIV, clock, 
            data_result, data_exception, data_resultRDY); 

    input [31:0] data_operandA, data_operandB;
    input ctrl_DIV, clock;

    output [31:0] data_result;
    output data_exception, data_resultRDY;

    


endmodule